module Program_Counter ();

endmodule
