/*
 * @file src/core/immext.v
 * @author Artin Zarei/Mohsen Mirzaei
 * @brief signed and unsigned extension.
 */

module ImmExt (
  input wire [15:0] immediate
);

  

endmodule
